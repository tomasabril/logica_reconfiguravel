library verilog;
use verilog.vl_types.all;
entity ex_1_logica_vlg_check_tst is
    port(
        AND_OUT         : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end ex_1_logica_vlg_check_tst;
