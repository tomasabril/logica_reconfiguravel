library verilog;
use verilog.vl_types.all;
entity ex_1_logica_vlg_vec_tst is
end ex_1_logica_vlg_vec_tst;
